// mysystem.v

// Generated using ACDS version 13.1 162 at 2015.01.22.17:35:24

`timescale 1 ps / 1 ps
module mysystem (
		input  wire        system_ref_clk_clk,      //    system_ref_clk.clk
		input  wire        system_ref_reset_reset,  //  system_ref_reset.reset
		output wire        sdram_clk_clk,           //         sdram_clk.clk
		output wire [12:0] memory_mem_a,            //            memory.mem_a
		output wire [2:0]  memory_mem_ba,           //                  .mem_ba
		output wire        memory_mem_ck,           //                  .mem_ck
		output wire        memory_mem_ck_n,         //                  .mem_ck_n
		output wire        memory_mem_cke,          //                  .mem_cke
		output wire        memory_mem_cs_n,         //                  .mem_cs_n
		output wire        memory_mem_ras_n,        //                  .mem_ras_n
		output wire        memory_mem_cas_n,        //                  .mem_cas_n
		output wire        memory_mem_we_n,         //                  .mem_we_n
		output wire        memory_mem_reset_n,      //                  .mem_reset_n
		inout  wire [7:0]  memory_mem_dq,           //                  .mem_dq
		inout  wire        memory_mem_dqs,          //                  .mem_dqs
		inout  wire        memory_mem_dqs_n,        //                  .mem_dqs_n
		output wire        memory_mem_odt,          //                  .mem_odt
		output wire        memory_mem_dm,           //                  .mem_dm
		input  wire        memory_oct_rzqin,        //                  .oct_rzqin
		input  wire        vga_pll_ref_clk_clk,     //   vga_pll_ref_clk.clk
		input  wire        vga_pll_ref_reset_reset, // vga_pll_ref_reset.reset
		output wire        vga_CLK,                 //               vga.CLK
		output wire        vga_HS,                  //                  .HS
		output wire        vga_VS,                  //                  .VS
		output wire        vga_BLANK,               //                  .BLANK
		output wire        vga_SYNC,                //                  .SYNC
		output wire [7:0]  vga_R,                   //                  .R
		output wire [7:0]  vga_G,                   //                  .G
		output wire [7:0]  vga_B,                   //                  .B
		output wire [12:0] sdram_addr,              //             sdram.addr
		output wire [1:0]  sdram_ba,                //                  .ba
		output wire        sdram_cas_n,             //                  .cas_n
		output wire        sdram_cke,               //                  .cke
		output wire        sdram_cs_n,              //                  .cs_n
		inout  wire [15:0] sdram_dq,                //                  .dq
		output wire [1:0]  sdram_dqm,               //                  .dqm
		output wire        sdram_ras_n,             //                  .ras_n
		output wire        sdram_we_n               //                  .we_n
	);

	wire          system_pll_sys_clk_clk;                                             // system_pll:sys_clk_clk -> [Onchip_SRAM:clk, Onchip_SRAM:clk2, SDRAM:clk, arm_a9_hps:f2h_axi_clk, arm_a9_hps:h2f_axi_clk, arm_a9_hps:h2f_lw_axi_clk, jtag_uart:clk, mm_interconnect_0:system_pll_sys_clk_clk, mm_interconnect_1:system_pll_sys_clk_clk, rst_controller:clk, rst_controller_002:clk, vgasystem_0:sys_clk_clk]
	wire          mm_interconnect_0_sdram_s1_waitrequest;                             // SDRAM:za_waitrequest -> mm_interconnect_0:SDRAM_s1_waitrequest
	wire   [15:0] mm_interconnect_0_sdram_s1_writedata;                               // mm_interconnect_0:SDRAM_s1_writedata -> SDRAM:az_data
	wire   [24:0] mm_interconnect_0_sdram_s1_address;                                 // mm_interconnect_0:SDRAM_s1_address -> SDRAM:az_addr
	wire          mm_interconnect_0_sdram_s1_chipselect;                              // mm_interconnect_0:SDRAM_s1_chipselect -> SDRAM:az_cs
	wire          mm_interconnect_0_sdram_s1_write;                                   // mm_interconnect_0:SDRAM_s1_write -> SDRAM:az_wr_n
	wire          mm_interconnect_0_sdram_s1_read;                                    // mm_interconnect_0:SDRAM_s1_read -> SDRAM:az_rd_n
	wire   [15:0] mm_interconnect_0_sdram_s1_readdata;                                // SDRAM:za_data -> mm_interconnect_0:SDRAM_s1_readdata
	wire          mm_interconnect_0_sdram_s1_readdatavalid;                           // SDRAM:za_valid -> mm_interconnect_0:SDRAM_s1_readdatavalid
	wire    [1:0] mm_interconnect_0_sdram_s1_byteenable;                              // mm_interconnect_0:SDRAM_s1_byteenable -> SDRAM:az_be_n
	wire          arm_a9_hps_h2f_axi_master_awvalid;                                  // arm_a9_hps:h2f_AWVALID -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_awvalid
	wire    [2:0] arm_a9_hps_h2f_axi_master_arsize;                                   // arm_a9_hps:h2f_ARSIZE -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_arsize
	wire    [1:0] arm_a9_hps_h2f_axi_master_arlock;                                   // arm_a9_hps:h2f_ARLOCK -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_arlock
	wire    [3:0] arm_a9_hps_h2f_axi_master_awcache;                                  // arm_a9_hps:h2f_AWCACHE -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_awcache
	wire          arm_a9_hps_h2f_axi_master_arready;                                  // mm_interconnect_0:arm_a9_hps_h2f_axi_master_arready -> arm_a9_hps:h2f_ARREADY
	wire   [11:0] arm_a9_hps_h2f_axi_master_arid;                                     // arm_a9_hps:h2f_ARID -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_arid
	wire          arm_a9_hps_h2f_axi_master_rready;                                   // arm_a9_hps:h2f_RREADY -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_rready
	wire          arm_a9_hps_h2f_axi_master_bready;                                   // arm_a9_hps:h2f_BREADY -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_bready
	wire    [2:0] arm_a9_hps_h2f_axi_master_awsize;                                   // arm_a9_hps:h2f_AWSIZE -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_awsize
	wire    [2:0] arm_a9_hps_h2f_axi_master_awprot;                                   // arm_a9_hps:h2f_AWPROT -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_awprot
	wire          arm_a9_hps_h2f_axi_master_arvalid;                                  // arm_a9_hps:h2f_ARVALID -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_arvalid
	wire    [2:0] arm_a9_hps_h2f_axi_master_arprot;                                   // arm_a9_hps:h2f_ARPROT -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_arprot
	wire   [11:0] arm_a9_hps_h2f_axi_master_bid;                                      // mm_interconnect_0:arm_a9_hps_h2f_axi_master_bid -> arm_a9_hps:h2f_BID
	wire    [3:0] arm_a9_hps_h2f_axi_master_arlen;                                    // arm_a9_hps:h2f_ARLEN -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_arlen
	wire          arm_a9_hps_h2f_axi_master_awready;                                  // mm_interconnect_0:arm_a9_hps_h2f_axi_master_awready -> arm_a9_hps:h2f_AWREADY
	wire   [11:0] arm_a9_hps_h2f_axi_master_awid;                                     // arm_a9_hps:h2f_AWID -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_awid
	wire          arm_a9_hps_h2f_axi_master_bvalid;                                   // mm_interconnect_0:arm_a9_hps_h2f_axi_master_bvalid -> arm_a9_hps:h2f_BVALID
	wire   [11:0] arm_a9_hps_h2f_axi_master_wid;                                      // arm_a9_hps:h2f_WID -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_wid
	wire    [1:0] arm_a9_hps_h2f_axi_master_awlock;                                   // arm_a9_hps:h2f_AWLOCK -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_awlock
	wire    [1:0] arm_a9_hps_h2f_axi_master_awburst;                                  // arm_a9_hps:h2f_AWBURST -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_awburst
	wire    [1:0] arm_a9_hps_h2f_axi_master_bresp;                                    // mm_interconnect_0:arm_a9_hps_h2f_axi_master_bresp -> arm_a9_hps:h2f_BRESP
	wire   [15:0] arm_a9_hps_h2f_axi_master_wstrb;                                    // arm_a9_hps:h2f_WSTRB -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_wstrb
	wire          arm_a9_hps_h2f_axi_master_rvalid;                                   // mm_interconnect_0:arm_a9_hps_h2f_axi_master_rvalid -> arm_a9_hps:h2f_RVALID
	wire  [127:0] arm_a9_hps_h2f_axi_master_wdata;                                    // arm_a9_hps:h2f_WDATA -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_wdata
	wire          arm_a9_hps_h2f_axi_master_wready;                                   // mm_interconnect_0:arm_a9_hps_h2f_axi_master_wready -> arm_a9_hps:h2f_WREADY
	wire    [1:0] arm_a9_hps_h2f_axi_master_arburst;                                  // arm_a9_hps:h2f_ARBURST -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_arburst
	wire  [127:0] arm_a9_hps_h2f_axi_master_rdata;                                    // mm_interconnect_0:arm_a9_hps_h2f_axi_master_rdata -> arm_a9_hps:h2f_RDATA
	wire   [29:0] arm_a9_hps_h2f_axi_master_araddr;                                   // arm_a9_hps:h2f_ARADDR -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_araddr
	wire    [3:0] arm_a9_hps_h2f_axi_master_arcache;                                  // arm_a9_hps:h2f_ARCACHE -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_arcache
	wire    [3:0] arm_a9_hps_h2f_axi_master_awlen;                                    // arm_a9_hps:h2f_AWLEN -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_awlen
	wire   [29:0] arm_a9_hps_h2f_axi_master_awaddr;                                   // arm_a9_hps:h2f_AWADDR -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_awaddr
	wire   [11:0] arm_a9_hps_h2f_axi_master_rid;                                      // mm_interconnect_0:arm_a9_hps_h2f_axi_master_rid -> arm_a9_hps:h2f_RID
	wire          arm_a9_hps_h2f_axi_master_wvalid;                                   // arm_a9_hps:h2f_WVALID -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_wvalid
	wire    [1:0] arm_a9_hps_h2f_axi_master_rresp;                                    // mm_interconnect_0:arm_a9_hps_h2f_axi_master_rresp -> arm_a9_hps:h2f_RRESP
	wire          arm_a9_hps_h2f_axi_master_wlast;                                    // arm_a9_hps:h2f_WLAST -> mm_interconnect_0:arm_a9_hps_h2f_axi_master_wlast
	wire          arm_a9_hps_h2f_axi_master_rlast;                                    // mm_interconnect_0:arm_a9_hps_h2f_axi_master_rlast -> arm_a9_hps:h2f_RLAST
	wire          vgasystem_0_pixel_dma_master_waitrequest;                           // mm_interconnect_0:vgasystem_0_pixel_dma_master_waitrequest -> vgasystem_0:pixel_dma_master_waitrequest
	wire   [31:0] vgasystem_0_pixel_dma_master_address;                               // vgasystem_0:pixel_dma_master_address -> mm_interconnect_0:vgasystem_0_pixel_dma_master_address
	wire          vgasystem_0_pixel_dma_master_lock;                                  // vgasystem_0:pixel_dma_master_lock -> mm_interconnect_0:vgasystem_0_pixel_dma_master_lock
	wire          vgasystem_0_pixel_dma_master_read;                                  // vgasystem_0:pixel_dma_master_read -> mm_interconnect_0:vgasystem_0_pixel_dma_master_read
	wire   [15:0] vgasystem_0_pixel_dma_master_readdata;                              // mm_interconnect_0:vgasystem_0_pixel_dma_master_readdata -> vgasystem_0:pixel_dma_master_readdata
	wire          vgasystem_0_pixel_dma_master_readdatavalid;                         // mm_interconnect_0:vgasystem_0_pixel_dma_master_readdatavalid -> vgasystem_0:pixel_dma_master_readdatavalid
	wire          mm_interconnect_0_vgasystem_0_char_buffer_slave_waitrequest;        // vgasystem_0:char_buffer_slave_waitrequest -> mm_interconnect_0:vgasystem_0_char_buffer_slave_waitrequest
	wire    [7:0] mm_interconnect_0_vgasystem_0_char_buffer_slave_writedata;          // mm_interconnect_0:vgasystem_0_char_buffer_slave_writedata -> vgasystem_0:char_buffer_slave_writedata
	wire   [12:0] mm_interconnect_0_vgasystem_0_char_buffer_slave_address;            // mm_interconnect_0:vgasystem_0_char_buffer_slave_address -> vgasystem_0:char_buffer_slave_address
	wire          mm_interconnect_0_vgasystem_0_char_buffer_slave_chipselect;         // mm_interconnect_0:vgasystem_0_char_buffer_slave_chipselect -> vgasystem_0:char_buffer_slave_chipselect
	wire          mm_interconnect_0_vgasystem_0_char_buffer_slave_write;              // mm_interconnect_0:vgasystem_0_char_buffer_slave_write -> vgasystem_0:char_buffer_slave_write
	wire          mm_interconnect_0_vgasystem_0_char_buffer_slave_read;               // mm_interconnect_0:vgasystem_0_char_buffer_slave_read -> vgasystem_0:char_buffer_slave_read
	wire    [7:0] mm_interconnect_0_vgasystem_0_char_buffer_slave_readdata;           // vgasystem_0:char_buffer_slave_readdata -> mm_interconnect_0:vgasystem_0_char_buffer_slave_readdata
	wire    [0:0] mm_interconnect_0_vgasystem_0_char_buffer_slave_byteenable;         // mm_interconnect_0:vgasystem_0_char_buffer_slave_byteenable -> vgasystem_0:char_buffer_slave_byteenable
	wire   [31:0] mm_interconnect_0_onchip_sram_s2_writedata;                         // mm_interconnect_0:Onchip_SRAM_s2_writedata -> Onchip_SRAM:writedata2
	wire   [11:0] mm_interconnect_0_onchip_sram_s2_address;                           // mm_interconnect_0:Onchip_SRAM_s2_address -> Onchip_SRAM:address2
	wire          mm_interconnect_0_onchip_sram_s2_chipselect;                        // mm_interconnect_0:Onchip_SRAM_s2_chipselect -> Onchip_SRAM:chipselect2
	wire          mm_interconnect_0_onchip_sram_s2_clken;                             // mm_interconnect_0:Onchip_SRAM_s2_clken -> Onchip_SRAM:clken2
	wire          mm_interconnect_0_onchip_sram_s2_write;                             // mm_interconnect_0:Onchip_SRAM_s2_write -> Onchip_SRAM:write2
	wire   [31:0] mm_interconnect_0_onchip_sram_s2_readdata;                          // Onchip_SRAM:readdata2 -> mm_interconnect_0:Onchip_SRAM_s2_readdata
	wire    [3:0] mm_interconnect_0_onchip_sram_s2_byteenable;                        // mm_interconnect_0:Onchip_SRAM_s2_byteenable -> Onchip_SRAM:byteenable2
	wire   [31:0] mm_interconnect_0_onchip_sram_s1_writedata;                         // mm_interconnect_0:Onchip_SRAM_s1_writedata -> Onchip_SRAM:writedata
	wire   [11:0] mm_interconnect_0_onchip_sram_s1_address;                           // mm_interconnect_0:Onchip_SRAM_s1_address -> Onchip_SRAM:address
	wire          mm_interconnect_0_onchip_sram_s1_chipselect;                        // mm_interconnect_0:Onchip_SRAM_s1_chipselect -> Onchip_SRAM:chipselect
	wire          mm_interconnect_0_onchip_sram_s1_clken;                             // mm_interconnect_0:Onchip_SRAM_s1_clken -> Onchip_SRAM:clken
	wire          mm_interconnect_0_onchip_sram_s1_write;                             // mm_interconnect_0:Onchip_SRAM_s1_write -> Onchip_SRAM:write
	wire   [31:0] mm_interconnect_0_onchip_sram_s1_readdata;                          // Onchip_SRAM:readdata -> mm_interconnect_0:Onchip_SRAM_s1_readdata
	wire    [3:0] mm_interconnect_0_onchip_sram_s1_byteenable;                        // mm_interconnect_0:Onchip_SRAM_s1_byteenable -> Onchip_SRAM:byteenable
	wire   [31:0] mm_interconnect_1_vgasystem_0_char_buffer_control_slave_writedata;  // mm_interconnect_1:vgasystem_0_char_buffer_control_slave_writedata -> vgasystem_0:char_buffer_control_slave_writedata
	wire    [0:0] mm_interconnect_1_vgasystem_0_char_buffer_control_slave_address;    // mm_interconnect_1:vgasystem_0_char_buffer_control_slave_address -> vgasystem_0:char_buffer_control_slave_address
	wire          mm_interconnect_1_vgasystem_0_char_buffer_control_slave_chipselect; // mm_interconnect_1:vgasystem_0_char_buffer_control_slave_chipselect -> vgasystem_0:char_buffer_control_slave_chipselect
	wire          mm_interconnect_1_vgasystem_0_char_buffer_control_slave_write;      // mm_interconnect_1:vgasystem_0_char_buffer_control_slave_write -> vgasystem_0:char_buffer_control_slave_write
	wire          mm_interconnect_1_vgasystem_0_char_buffer_control_slave_read;       // mm_interconnect_1:vgasystem_0_char_buffer_control_slave_read -> vgasystem_0:char_buffer_control_slave_read
	wire   [31:0] mm_interconnect_1_vgasystem_0_char_buffer_control_slave_readdata;   // vgasystem_0:char_buffer_control_slave_readdata -> mm_interconnect_1:vgasystem_0_char_buffer_control_slave_readdata
	wire    [3:0] mm_interconnect_1_vgasystem_0_char_buffer_control_slave_byteenable; // mm_interconnect_1:vgasystem_0_char_buffer_control_slave_byteenable -> vgasystem_0:char_buffer_control_slave_byteenable
	wire   [31:0] mm_interconnect_1_vgasystem_0_pixel_dma_control_slave_writedata;    // mm_interconnect_1:vgasystem_0_pixel_dma_control_slave_writedata -> vgasystem_0:pixel_dma_control_slave_writedata
	wire    [1:0] mm_interconnect_1_vgasystem_0_pixel_dma_control_slave_address;      // mm_interconnect_1:vgasystem_0_pixel_dma_control_slave_address -> vgasystem_0:pixel_dma_control_slave_address
	wire          mm_interconnect_1_vgasystem_0_pixel_dma_control_slave_write;        // mm_interconnect_1:vgasystem_0_pixel_dma_control_slave_write -> vgasystem_0:pixel_dma_control_slave_write
	wire          mm_interconnect_1_vgasystem_0_pixel_dma_control_slave_read;         // mm_interconnect_1:vgasystem_0_pixel_dma_control_slave_read -> vgasystem_0:pixel_dma_control_slave_read
	wire   [31:0] mm_interconnect_1_vgasystem_0_pixel_dma_control_slave_readdata;     // vgasystem_0:pixel_dma_control_slave_readdata -> mm_interconnect_1:vgasystem_0_pixel_dma_control_slave_readdata
	wire    [3:0] mm_interconnect_1_vgasystem_0_pixel_dma_control_slave_byteenable;   // mm_interconnect_1:vgasystem_0_pixel_dma_control_slave_byteenable -> vgasystem_0:pixel_dma_control_slave_byteenable
	wire          arm_a9_hps_h2f_lw_axi_master_awvalid;                               // arm_a9_hps:h2f_lw_AWVALID -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_awvalid
	wire    [2:0] arm_a9_hps_h2f_lw_axi_master_arsize;                                // arm_a9_hps:h2f_lw_ARSIZE -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_arsize
	wire    [1:0] arm_a9_hps_h2f_lw_axi_master_arlock;                                // arm_a9_hps:h2f_lw_ARLOCK -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_arlock
	wire    [3:0] arm_a9_hps_h2f_lw_axi_master_awcache;                               // arm_a9_hps:h2f_lw_AWCACHE -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_awcache
	wire          arm_a9_hps_h2f_lw_axi_master_arready;                               // mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_arready -> arm_a9_hps:h2f_lw_ARREADY
	wire   [11:0] arm_a9_hps_h2f_lw_axi_master_arid;                                  // arm_a9_hps:h2f_lw_ARID -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_arid
	wire          arm_a9_hps_h2f_lw_axi_master_rready;                                // arm_a9_hps:h2f_lw_RREADY -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_rready
	wire          arm_a9_hps_h2f_lw_axi_master_bready;                                // arm_a9_hps:h2f_lw_BREADY -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_bready
	wire    [2:0] arm_a9_hps_h2f_lw_axi_master_awsize;                                // arm_a9_hps:h2f_lw_AWSIZE -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_awsize
	wire    [2:0] arm_a9_hps_h2f_lw_axi_master_awprot;                                // arm_a9_hps:h2f_lw_AWPROT -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_awprot
	wire          arm_a9_hps_h2f_lw_axi_master_arvalid;                               // arm_a9_hps:h2f_lw_ARVALID -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_arvalid
	wire    [2:0] arm_a9_hps_h2f_lw_axi_master_arprot;                                // arm_a9_hps:h2f_lw_ARPROT -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_arprot
	wire   [11:0] arm_a9_hps_h2f_lw_axi_master_bid;                                   // mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_bid -> arm_a9_hps:h2f_lw_BID
	wire    [3:0] arm_a9_hps_h2f_lw_axi_master_arlen;                                 // arm_a9_hps:h2f_lw_ARLEN -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_arlen
	wire          arm_a9_hps_h2f_lw_axi_master_awready;                               // mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_awready -> arm_a9_hps:h2f_lw_AWREADY
	wire   [11:0] arm_a9_hps_h2f_lw_axi_master_awid;                                  // arm_a9_hps:h2f_lw_AWID -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_awid
	wire          arm_a9_hps_h2f_lw_axi_master_bvalid;                                // mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_bvalid -> arm_a9_hps:h2f_lw_BVALID
	wire   [11:0] arm_a9_hps_h2f_lw_axi_master_wid;                                   // arm_a9_hps:h2f_lw_WID -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_wid
	wire    [1:0] arm_a9_hps_h2f_lw_axi_master_awlock;                                // arm_a9_hps:h2f_lw_AWLOCK -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_awlock
	wire    [1:0] arm_a9_hps_h2f_lw_axi_master_awburst;                               // arm_a9_hps:h2f_lw_AWBURST -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_awburst
	wire    [1:0] arm_a9_hps_h2f_lw_axi_master_bresp;                                 // mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_bresp -> arm_a9_hps:h2f_lw_BRESP
	wire    [3:0] arm_a9_hps_h2f_lw_axi_master_wstrb;                                 // arm_a9_hps:h2f_lw_WSTRB -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_wstrb
	wire          arm_a9_hps_h2f_lw_axi_master_rvalid;                                // mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_rvalid -> arm_a9_hps:h2f_lw_RVALID
	wire   [31:0] arm_a9_hps_h2f_lw_axi_master_wdata;                                 // arm_a9_hps:h2f_lw_WDATA -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_wdata
	wire          arm_a9_hps_h2f_lw_axi_master_wready;                                // mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_wready -> arm_a9_hps:h2f_lw_WREADY
	wire    [1:0] arm_a9_hps_h2f_lw_axi_master_arburst;                               // arm_a9_hps:h2f_lw_ARBURST -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_arburst
	wire   [31:0] arm_a9_hps_h2f_lw_axi_master_rdata;                                 // mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_rdata -> arm_a9_hps:h2f_lw_RDATA
	wire   [20:0] arm_a9_hps_h2f_lw_axi_master_araddr;                                // arm_a9_hps:h2f_lw_ARADDR -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_araddr
	wire    [3:0] arm_a9_hps_h2f_lw_axi_master_arcache;                               // arm_a9_hps:h2f_lw_ARCACHE -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_arcache
	wire    [3:0] arm_a9_hps_h2f_lw_axi_master_awlen;                                 // arm_a9_hps:h2f_lw_AWLEN -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_awlen
	wire   [20:0] arm_a9_hps_h2f_lw_axi_master_awaddr;                                // arm_a9_hps:h2f_lw_AWADDR -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_awaddr
	wire   [11:0] arm_a9_hps_h2f_lw_axi_master_rid;                                   // mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_rid -> arm_a9_hps:h2f_lw_RID
	wire          arm_a9_hps_h2f_lw_axi_master_wvalid;                                // arm_a9_hps:h2f_lw_WVALID -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_wvalid
	wire    [1:0] arm_a9_hps_h2f_lw_axi_master_rresp;                                 // mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_rresp -> arm_a9_hps:h2f_lw_RRESP
	wire          arm_a9_hps_h2f_lw_axi_master_wlast;                                 // arm_a9_hps:h2f_lw_WLAST -> mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_wlast
	wire          arm_a9_hps_h2f_lw_axi_master_rlast;                                 // mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_rlast -> arm_a9_hps:h2f_lw_RLAST
	wire          mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest;          // jtag_uart:av_waitrequest -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata;            // mm_interconnect_1:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire    [0:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_address;              // mm_interconnect_1:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire          mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect;           // mm_interconnect_1:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire          mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;                // mm_interconnect_1:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire          mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;                 // mm_interconnect_1:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire   [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata;             // jtag_uart:av_readdata -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_readdata
	wire          irq_mapper_receiver0_irq;                                           // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire   [31:0] arm_a9_hps_f2h_irq0_irq;                                            // irq_mapper:sender_irq -> arm_a9_hps:f2h_irq_p0
	wire   [31:0] arm_a9_hps_f2h_irq1_irq;                                            // irq_mapper_001:sender_irq -> arm_a9_hps:f2h_irq_p1
	wire          rst_controller_reset_out_reset;                                     // rst_controller:reset_out -> [Onchip_SRAM:reset, Onchip_SRAM:reset2, SDRAM:reset_n, jtag_uart:rst_n, mm_interconnect_0:Onchip_SRAM_reset1_reset_bridge_in_reset_reset, mm_interconnect_0:vgasystem_0_sys_reset_reset_bridge_in_reset_reset, mm_interconnect_1:jtag_uart_reset_reset_bridge_in_reset_reset, mm_interconnect_1:vgasystem_0_sys_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire          rst_controller_reset_out_reset_req;                                 // rst_controller:reset_req -> [Onchip_SRAM:reset_req, Onchip_SRAM:reset_req2, rst_translator:reset_req_in]
	wire          system_pll_reset_source_reset;                                      // system_pll:reset_source_reset -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	wire          arm_a9_hps_h2f_reset_reset;                                         // arm_a9_hps:h2f_rst_n -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in0]
	wire          rst_controller_001_reset_out_reset;                                 // rst_controller_001:reset_out -> vgasystem_0:sys_reset_reset_n
	wire          rst_controller_002_reset_out_reset;                                 // rst_controller_002:reset_out -> [mm_interconnect_0:arm_a9_hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:arm_a9_hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]

	mysystem_system_pll system_pll (
		.ref_clk_clk        (system_ref_clk_clk),            //      ref_clk.clk
		.ref_reset_reset    (system_ref_reset_reset),        //    ref_reset.reset
		.sys_clk_clk        (system_pll_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),                 //    sdram_clk.clk
		.reset_source_reset (system_pll_reset_source_reset)  // reset_source.reset
	);

	mysystem_arm_a9_hps #(
		.F2S_Width (2),
		.S2F_Width (3)
	) arm_a9_hps (
		.mem_a          (memory_mem_a),                         //            memory.mem_a
		.mem_ba         (memory_mem_ba),                        //                  .mem_ba
		.mem_ck         (memory_mem_ck),                        //                  .mem_ck
		.mem_ck_n       (memory_mem_ck_n),                      //                  .mem_ck_n
		.mem_cke        (memory_mem_cke),                       //                  .mem_cke
		.mem_cs_n       (memory_mem_cs_n),                      //                  .mem_cs_n
		.mem_ras_n      (memory_mem_ras_n),                     //                  .mem_ras_n
		.mem_cas_n      (memory_mem_cas_n),                     //                  .mem_cas_n
		.mem_we_n       (memory_mem_we_n),                      //                  .mem_we_n
		.mem_reset_n    (memory_mem_reset_n),                   //                  .mem_reset_n
		.mem_dq         (memory_mem_dq),                        //                  .mem_dq
		.mem_dqs        (memory_mem_dqs),                       //                  .mem_dqs
		.mem_dqs_n      (memory_mem_dqs_n),                     //                  .mem_dqs_n
		.mem_odt        (memory_mem_odt),                       //                  .mem_odt
		.mem_dm         (memory_mem_dm),                        //                  .mem_dm
		.oct_rzqin      (memory_oct_rzqin),                     //                  .oct_rzqin
		.h2f_rst_n      (arm_a9_hps_h2f_reset_reset),           //         h2f_reset.reset_n
		.h2f_axi_clk    (system_pll_sys_clk_clk),               //     h2f_axi_clock.clk
		.h2f_AWID       (arm_a9_hps_h2f_axi_master_awid),       //    h2f_axi_master.awid
		.h2f_AWADDR     (arm_a9_hps_h2f_axi_master_awaddr),     //                  .awaddr
		.h2f_AWLEN      (arm_a9_hps_h2f_axi_master_awlen),      //                  .awlen
		.h2f_AWSIZE     (arm_a9_hps_h2f_axi_master_awsize),     //                  .awsize
		.h2f_AWBURST    (arm_a9_hps_h2f_axi_master_awburst),    //                  .awburst
		.h2f_AWLOCK     (arm_a9_hps_h2f_axi_master_awlock),     //                  .awlock
		.h2f_AWCACHE    (arm_a9_hps_h2f_axi_master_awcache),    //                  .awcache
		.h2f_AWPROT     (arm_a9_hps_h2f_axi_master_awprot),     //                  .awprot
		.h2f_AWVALID    (arm_a9_hps_h2f_axi_master_awvalid),    //                  .awvalid
		.h2f_AWREADY    (arm_a9_hps_h2f_axi_master_awready),    //                  .awready
		.h2f_WID        (arm_a9_hps_h2f_axi_master_wid),        //                  .wid
		.h2f_WDATA      (arm_a9_hps_h2f_axi_master_wdata),      //                  .wdata
		.h2f_WSTRB      (arm_a9_hps_h2f_axi_master_wstrb),      //                  .wstrb
		.h2f_WLAST      (arm_a9_hps_h2f_axi_master_wlast),      //                  .wlast
		.h2f_WVALID     (arm_a9_hps_h2f_axi_master_wvalid),     //                  .wvalid
		.h2f_WREADY     (arm_a9_hps_h2f_axi_master_wready),     //                  .wready
		.h2f_BID        (arm_a9_hps_h2f_axi_master_bid),        //                  .bid
		.h2f_BRESP      (arm_a9_hps_h2f_axi_master_bresp),      //                  .bresp
		.h2f_BVALID     (arm_a9_hps_h2f_axi_master_bvalid),     //                  .bvalid
		.h2f_BREADY     (arm_a9_hps_h2f_axi_master_bready),     //                  .bready
		.h2f_ARID       (arm_a9_hps_h2f_axi_master_arid),       //                  .arid
		.h2f_ARADDR     (arm_a9_hps_h2f_axi_master_araddr),     //                  .araddr
		.h2f_ARLEN      (arm_a9_hps_h2f_axi_master_arlen),      //                  .arlen
		.h2f_ARSIZE     (arm_a9_hps_h2f_axi_master_arsize),     //                  .arsize
		.h2f_ARBURST    (arm_a9_hps_h2f_axi_master_arburst),    //                  .arburst
		.h2f_ARLOCK     (arm_a9_hps_h2f_axi_master_arlock),     //                  .arlock
		.h2f_ARCACHE    (arm_a9_hps_h2f_axi_master_arcache),    //                  .arcache
		.h2f_ARPROT     (arm_a9_hps_h2f_axi_master_arprot),     //                  .arprot
		.h2f_ARVALID    (arm_a9_hps_h2f_axi_master_arvalid),    //                  .arvalid
		.h2f_ARREADY    (arm_a9_hps_h2f_axi_master_arready),    //                  .arready
		.h2f_RID        (arm_a9_hps_h2f_axi_master_rid),        //                  .rid
		.h2f_RDATA      (arm_a9_hps_h2f_axi_master_rdata),      //                  .rdata
		.h2f_RRESP      (arm_a9_hps_h2f_axi_master_rresp),      //                  .rresp
		.h2f_RLAST      (arm_a9_hps_h2f_axi_master_rlast),      //                  .rlast
		.h2f_RVALID     (arm_a9_hps_h2f_axi_master_rvalid),     //                  .rvalid
		.h2f_RREADY     (arm_a9_hps_h2f_axi_master_rready),     //                  .rready
		.f2h_axi_clk    (system_pll_sys_clk_clk),               //     f2h_axi_clock.clk
		.f2h_AWID       (),                                     //     f2h_axi_slave.awid
		.f2h_AWADDR     (),                                     //                  .awaddr
		.f2h_AWLEN      (),                                     //                  .awlen
		.f2h_AWSIZE     (),                                     //                  .awsize
		.f2h_AWBURST    (),                                     //                  .awburst
		.f2h_AWLOCK     (),                                     //                  .awlock
		.f2h_AWCACHE    (),                                     //                  .awcache
		.f2h_AWPROT     (),                                     //                  .awprot
		.f2h_AWVALID    (),                                     //                  .awvalid
		.f2h_AWREADY    (),                                     //                  .awready
		.f2h_AWUSER     (),                                     //                  .awuser
		.f2h_WID        (),                                     //                  .wid
		.f2h_WDATA      (),                                     //                  .wdata
		.f2h_WSTRB      (),                                     //                  .wstrb
		.f2h_WLAST      (),                                     //                  .wlast
		.f2h_WVALID     (),                                     //                  .wvalid
		.f2h_WREADY     (),                                     //                  .wready
		.f2h_BID        (),                                     //                  .bid
		.f2h_BRESP      (),                                     //                  .bresp
		.f2h_BVALID     (),                                     //                  .bvalid
		.f2h_BREADY     (),                                     //                  .bready
		.f2h_ARID       (),                                     //                  .arid
		.f2h_ARADDR     (),                                     //                  .araddr
		.f2h_ARLEN      (),                                     //                  .arlen
		.f2h_ARSIZE     (),                                     //                  .arsize
		.f2h_ARBURST    (),                                     //                  .arburst
		.f2h_ARLOCK     (),                                     //                  .arlock
		.f2h_ARCACHE    (),                                     //                  .arcache
		.f2h_ARPROT     (),                                     //                  .arprot
		.f2h_ARVALID    (),                                     //                  .arvalid
		.f2h_ARREADY    (),                                     //                  .arready
		.f2h_ARUSER     (),                                     //                  .aruser
		.f2h_RID        (),                                     //                  .rid
		.f2h_RDATA      (),                                     //                  .rdata
		.f2h_RRESP      (),                                     //                  .rresp
		.f2h_RLAST      (),                                     //                  .rlast
		.f2h_RVALID     (),                                     //                  .rvalid
		.f2h_RREADY     (),                                     //                  .rready
		.h2f_lw_axi_clk (system_pll_sys_clk_clk),               //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID    (arm_a9_hps_h2f_lw_axi_master_awid),    // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR  (arm_a9_hps_h2f_lw_axi_master_awaddr),  //                  .awaddr
		.h2f_lw_AWLEN   (arm_a9_hps_h2f_lw_axi_master_awlen),   //                  .awlen
		.h2f_lw_AWSIZE  (arm_a9_hps_h2f_lw_axi_master_awsize),  //                  .awsize
		.h2f_lw_AWBURST (arm_a9_hps_h2f_lw_axi_master_awburst), //                  .awburst
		.h2f_lw_AWLOCK  (arm_a9_hps_h2f_lw_axi_master_awlock),  //                  .awlock
		.h2f_lw_AWCACHE (arm_a9_hps_h2f_lw_axi_master_awcache), //                  .awcache
		.h2f_lw_AWPROT  (arm_a9_hps_h2f_lw_axi_master_awprot),  //                  .awprot
		.h2f_lw_AWVALID (arm_a9_hps_h2f_lw_axi_master_awvalid), //                  .awvalid
		.h2f_lw_AWREADY (arm_a9_hps_h2f_lw_axi_master_awready), //                  .awready
		.h2f_lw_WID     (arm_a9_hps_h2f_lw_axi_master_wid),     //                  .wid
		.h2f_lw_WDATA   (arm_a9_hps_h2f_lw_axi_master_wdata),   //                  .wdata
		.h2f_lw_WSTRB   (arm_a9_hps_h2f_lw_axi_master_wstrb),   //                  .wstrb
		.h2f_lw_WLAST   (arm_a9_hps_h2f_lw_axi_master_wlast),   //                  .wlast
		.h2f_lw_WVALID  (arm_a9_hps_h2f_lw_axi_master_wvalid),  //                  .wvalid
		.h2f_lw_WREADY  (arm_a9_hps_h2f_lw_axi_master_wready),  //                  .wready
		.h2f_lw_BID     (arm_a9_hps_h2f_lw_axi_master_bid),     //                  .bid
		.h2f_lw_BRESP   (arm_a9_hps_h2f_lw_axi_master_bresp),   //                  .bresp
		.h2f_lw_BVALID  (arm_a9_hps_h2f_lw_axi_master_bvalid),  //                  .bvalid
		.h2f_lw_BREADY  (arm_a9_hps_h2f_lw_axi_master_bready),  //                  .bready
		.h2f_lw_ARID    (arm_a9_hps_h2f_lw_axi_master_arid),    //                  .arid
		.h2f_lw_ARADDR  (arm_a9_hps_h2f_lw_axi_master_araddr),  //                  .araddr
		.h2f_lw_ARLEN   (arm_a9_hps_h2f_lw_axi_master_arlen),   //                  .arlen
		.h2f_lw_ARSIZE  (arm_a9_hps_h2f_lw_axi_master_arsize),  //                  .arsize
		.h2f_lw_ARBURST (arm_a9_hps_h2f_lw_axi_master_arburst), //                  .arburst
		.h2f_lw_ARLOCK  (arm_a9_hps_h2f_lw_axi_master_arlock),  //                  .arlock
		.h2f_lw_ARCACHE (arm_a9_hps_h2f_lw_axi_master_arcache), //                  .arcache
		.h2f_lw_ARPROT  (arm_a9_hps_h2f_lw_axi_master_arprot),  //                  .arprot
		.h2f_lw_ARVALID (arm_a9_hps_h2f_lw_axi_master_arvalid), //                  .arvalid
		.h2f_lw_ARREADY (arm_a9_hps_h2f_lw_axi_master_arready), //                  .arready
		.h2f_lw_RID     (arm_a9_hps_h2f_lw_axi_master_rid),     //                  .rid
		.h2f_lw_RDATA   (arm_a9_hps_h2f_lw_axi_master_rdata),   //                  .rdata
		.h2f_lw_RRESP   (arm_a9_hps_h2f_lw_axi_master_rresp),   //                  .rresp
		.h2f_lw_RLAST   (arm_a9_hps_h2f_lw_axi_master_rlast),   //                  .rlast
		.h2f_lw_RVALID  (arm_a9_hps_h2f_lw_axi_master_rvalid),  //                  .rvalid
		.h2f_lw_RREADY  (arm_a9_hps_h2f_lw_axi_master_rready),  //                  .rready
		.f2h_irq_p0     (arm_a9_hps_f2h_irq0_irq),              //          f2h_irq0.irq
		.f2h_irq_p1     (arm_a9_hps_f2h_irq1_irq)               //          f2h_irq1.irq
	);

	mysystem_Onchip_SRAM onchip_sram (
		.clk         (system_pll_sys_clk_clk),                      //   clk1.clk
		.address     (mm_interconnect_0_onchip_sram_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_onchip_sram_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_onchip_sram_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_onchip_sram_s1_write),      //       .write
		.readdata    (mm_interconnect_0_onchip_sram_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_onchip_sram_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_onchip_sram_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),              // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),          //       .reset_req
		.address2    (mm_interconnect_0_onchip_sram_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_onchip_sram_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_onchip_sram_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_onchip_sram_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_onchip_sram_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_onchip_sram_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_onchip_sram_s2_byteenable), //       .byteenable
		.clk2        (system_pll_sys_clk_clk),                      //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),              // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req)           //       .reset_req
	);

	mysystem_jtag_uart jtag_uart (
		.clk            (system_pll_sys_clk_clk),                                    //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	mysystem_vgasystem_0 vgasystem_0 (
		.sys_clk_clk                          (system_pll_sys_clk_clk),                                             //                   sys_clk.clk
		.sys_reset_reset_n                    (~rst_controller_001_reset_out_reset),                                //                 sys_reset.reset_n
		.vga_pll_ref_clk_clk                  (vga_pll_ref_clk_clk),                                                //           vga_pll_ref_clk.clk
		.vga_pll_ref_reset_reset              (vga_pll_ref_reset_reset),                                            //         vga_pll_ref_reset.reset
		.pixel_dma_master_readdatavalid       (vgasystem_0_pixel_dma_master_readdatavalid),                         //          pixel_dma_master.readdatavalid
		.pixel_dma_master_waitrequest         (vgasystem_0_pixel_dma_master_waitrequest),                           //                          .waitrequest
		.pixel_dma_master_address             (vgasystem_0_pixel_dma_master_address),                               //                          .address
		.pixel_dma_master_lock                (vgasystem_0_pixel_dma_master_lock),                                  //                          .lock
		.pixel_dma_master_read                (vgasystem_0_pixel_dma_master_read),                                  //                          .read
		.pixel_dma_master_readdata            (vgasystem_0_pixel_dma_master_readdata),                              //                          .readdata
		.pixel_dma_control_slave_address      (mm_interconnect_1_vgasystem_0_pixel_dma_control_slave_address),      //   pixel_dma_control_slave.address
		.pixel_dma_control_slave_byteenable   (mm_interconnect_1_vgasystem_0_pixel_dma_control_slave_byteenable),   //                          .byteenable
		.pixel_dma_control_slave_read         (mm_interconnect_1_vgasystem_0_pixel_dma_control_slave_read),         //                          .read
		.pixel_dma_control_slave_write        (mm_interconnect_1_vgasystem_0_pixel_dma_control_slave_write),        //                          .write
		.pixel_dma_control_slave_writedata    (mm_interconnect_1_vgasystem_0_pixel_dma_control_slave_writedata),    //                          .writedata
		.pixel_dma_control_slave_readdata     (mm_interconnect_1_vgasystem_0_pixel_dma_control_slave_readdata),     //                          .readdata
		.char_buffer_control_slave_address    (mm_interconnect_1_vgasystem_0_char_buffer_control_slave_address),    // char_buffer_control_slave.address
		.char_buffer_control_slave_byteenable (mm_interconnect_1_vgasystem_0_char_buffer_control_slave_byteenable), //                          .byteenable
		.char_buffer_control_slave_chipselect (mm_interconnect_1_vgasystem_0_char_buffer_control_slave_chipselect), //                          .chipselect
		.char_buffer_control_slave_read       (mm_interconnect_1_vgasystem_0_char_buffer_control_slave_read),       //                          .read
		.char_buffer_control_slave_write      (mm_interconnect_1_vgasystem_0_char_buffer_control_slave_write),      //                          .write
		.char_buffer_control_slave_writedata  (mm_interconnect_1_vgasystem_0_char_buffer_control_slave_writedata),  //                          .writedata
		.char_buffer_control_slave_readdata   (mm_interconnect_1_vgasystem_0_char_buffer_control_slave_readdata),   //                          .readdata
		.char_buffer_slave_byteenable         (mm_interconnect_0_vgasystem_0_char_buffer_slave_byteenable),         //         char_buffer_slave.byteenable
		.char_buffer_slave_chipselect         (mm_interconnect_0_vgasystem_0_char_buffer_slave_chipselect),         //                          .chipselect
		.char_buffer_slave_read               (mm_interconnect_0_vgasystem_0_char_buffer_slave_read),               //                          .read
		.char_buffer_slave_write              (mm_interconnect_0_vgasystem_0_char_buffer_slave_write),              //                          .write
		.char_buffer_slave_writedata          (mm_interconnect_0_vgasystem_0_char_buffer_slave_writedata),          //                          .writedata
		.char_buffer_slave_readdata           (mm_interconnect_0_vgasystem_0_char_buffer_slave_readdata),           //                          .readdata
		.char_buffer_slave_waitrequest        (mm_interconnect_0_vgasystem_0_char_buffer_slave_waitrequest),        //                          .waitrequest
		.char_buffer_slave_address            (mm_interconnect_0_vgasystem_0_char_buffer_slave_address),            //                          .address
		.vga_CLK                              (vga_CLK),                                                            //                       vga.CLK
		.vga_HS                               (vga_HS),                                                             //                          .HS
		.vga_VS                               (vga_VS),                                                             //                          .VS
		.vga_BLANK                            (vga_BLANK),                                                          //                          .BLANK
		.vga_SYNC                             (vga_SYNC),                                                           //                          .SYNC
		.vga_R                                (vga_R),                                                              //                          .R
		.vga_G                                (vga_G),                                                              //                          .G
		.vga_B                                (vga_B)                                                               //                          .B
	);

	mysystem_SDRAM sdram (
		.clk            (system_pll_sys_clk_clk),                   //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	mysystem_mm_interconnect_0 mm_interconnect_0 (
		.arm_a9_hps_h2f_axi_master_awid                                        (arm_a9_hps_h2f_axi_master_awid),                              //                                       arm_a9_hps_h2f_axi_master.awid
		.arm_a9_hps_h2f_axi_master_awaddr                                      (arm_a9_hps_h2f_axi_master_awaddr),                            //                                                                .awaddr
		.arm_a9_hps_h2f_axi_master_awlen                                       (arm_a9_hps_h2f_axi_master_awlen),                             //                                                                .awlen
		.arm_a9_hps_h2f_axi_master_awsize                                      (arm_a9_hps_h2f_axi_master_awsize),                            //                                                                .awsize
		.arm_a9_hps_h2f_axi_master_awburst                                     (arm_a9_hps_h2f_axi_master_awburst),                           //                                                                .awburst
		.arm_a9_hps_h2f_axi_master_awlock                                      (arm_a9_hps_h2f_axi_master_awlock),                            //                                                                .awlock
		.arm_a9_hps_h2f_axi_master_awcache                                     (arm_a9_hps_h2f_axi_master_awcache),                           //                                                                .awcache
		.arm_a9_hps_h2f_axi_master_awprot                                      (arm_a9_hps_h2f_axi_master_awprot),                            //                                                                .awprot
		.arm_a9_hps_h2f_axi_master_awvalid                                     (arm_a9_hps_h2f_axi_master_awvalid),                           //                                                                .awvalid
		.arm_a9_hps_h2f_axi_master_awready                                     (arm_a9_hps_h2f_axi_master_awready),                           //                                                                .awready
		.arm_a9_hps_h2f_axi_master_wid                                         (arm_a9_hps_h2f_axi_master_wid),                               //                                                                .wid
		.arm_a9_hps_h2f_axi_master_wdata                                       (arm_a9_hps_h2f_axi_master_wdata),                             //                                                                .wdata
		.arm_a9_hps_h2f_axi_master_wstrb                                       (arm_a9_hps_h2f_axi_master_wstrb),                             //                                                                .wstrb
		.arm_a9_hps_h2f_axi_master_wlast                                       (arm_a9_hps_h2f_axi_master_wlast),                             //                                                                .wlast
		.arm_a9_hps_h2f_axi_master_wvalid                                      (arm_a9_hps_h2f_axi_master_wvalid),                            //                                                                .wvalid
		.arm_a9_hps_h2f_axi_master_wready                                      (arm_a9_hps_h2f_axi_master_wready),                            //                                                                .wready
		.arm_a9_hps_h2f_axi_master_bid                                         (arm_a9_hps_h2f_axi_master_bid),                               //                                                                .bid
		.arm_a9_hps_h2f_axi_master_bresp                                       (arm_a9_hps_h2f_axi_master_bresp),                             //                                                                .bresp
		.arm_a9_hps_h2f_axi_master_bvalid                                      (arm_a9_hps_h2f_axi_master_bvalid),                            //                                                                .bvalid
		.arm_a9_hps_h2f_axi_master_bready                                      (arm_a9_hps_h2f_axi_master_bready),                            //                                                                .bready
		.arm_a9_hps_h2f_axi_master_arid                                        (arm_a9_hps_h2f_axi_master_arid),                              //                                                                .arid
		.arm_a9_hps_h2f_axi_master_araddr                                      (arm_a9_hps_h2f_axi_master_araddr),                            //                                                                .araddr
		.arm_a9_hps_h2f_axi_master_arlen                                       (arm_a9_hps_h2f_axi_master_arlen),                             //                                                                .arlen
		.arm_a9_hps_h2f_axi_master_arsize                                      (arm_a9_hps_h2f_axi_master_arsize),                            //                                                                .arsize
		.arm_a9_hps_h2f_axi_master_arburst                                     (arm_a9_hps_h2f_axi_master_arburst),                           //                                                                .arburst
		.arm_a9_hps_h2f_axi_master_arlock                                      (arm_a9_hps_h2f_axi_master_arlock),                            //                                                                .arlock
		.arm_a9_hps_h2f_axi_master_arcache                                     (arm_a9_hps_h2f_axi_master_arcache),                           //                                                                .arcache
		.arm_a9_hps_h2f_axi_master_arprot                                      (arm_a9_hps_h2f_axi_master_arprot),                            //                                                                .arprot
		.arm_a9_hps_h2f_axi_master_arvalid                                     (arm_a9_hps_h2f_axi_master_arvalid),                           //                                                                .arvalid
		.arm_a9_hps_h2f_axi_master_arready                                     (arm_a9_hps_h2f_axi_master_arready),                           //                                                                .arready
		.arm_a9_hps_h2f_axi_master_rid                                         (arm_a9_hps_h2f_axi_master_rid),                               //                                                                .rid
		.arm_a9_hps_h2f_axi_master_rdata                                       (arm_a9_hps_h2f_axi_master_rdata),                             //                                                                .rdata
		.arm_a9_hps_h2f_axi_master_rresp                                       (arm_a9_hps_h2f_axi_master_rresp),                             //                                                                .rresp
		.arm_a9_hps_h2f_axi_master_rlast                                       (arm_a9_hps_h2f_axi_master_rlast),                             //                                                                .rlast
		.arm_a9_hps_h2f_axi_master_rvalid                                      (arm_a9_hps_h2f_axi_master_rvalid),                            //                                                                .rvalid
		.arm_a9_hps_h2f_axi_master_rready                                      (arm_a9_hps_h2f_axi_master_rready),                            //                                                                .rready
		.system_pll_sys_clk_clk                                                (system_pll_sys_clk_clk),                                      //                                              system_pll_sys_clk.clk
		.arm_a9_hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                          // arm_a9_hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.Onchip_SRAM_reset1_reset_bridge_in_reset_reset                        (rst_controller_reset_out_reset),                              //                        Onchip_SRAM_reset1_reset_bridge_in_reset.reset
		.vgasystem_0_sys_reset_reset_bridge_in_reset_reset                     (rst_controller_reset_out_reset),                              //                     vgasystem_0_sys_reset_reset_bridge_in_reset.reset
		.vgasystem_0_pixel_dma_master_address                                  (vgasystem_0_pixel_dma_master_address),                        //                                    vgasystem_0_pixel_dma_master.address
		.vgasystem_0_pixel_dma_master_waitrequest                              (vgasystem_0_pixel_dma_master_waitrequest),                    //                                                                .waitrequest
		.vgasystem_0_pixel_dma_master_read                                     (vgasystem_0_pixel_dma_master_read),                           //                                                                .read
		.vgasystem_0_pixel_dma_master_readdata                                 (vgasystem_0_pixel_dma_master_readdata),                       //                                                                .readdata
		.vgasystem_0_pixel_dma_master_readdatavalid                            (vgasystem_0_pixel_dma_master_readdatavalid),                  //                                                                .readdatavalid
		.vgasystem_0_pixel_dma_master_lock                                     (vgasystem_0_pixel_dma_master_lock),                           //                                                                .lock
		.Onchip_SRAM_s1_address                                                (mm_interconnect_0_onchip_sram_s1_address),                    //                                                  Onchip_SRAM_s1.address
		.Onchip_SRAM_s1_write                                                  (mm_interconnect_0_onchip_sram_s1_write),                      //                                                                .write
		.Onchip_SRAM_s1_readdata                                               (mm_interconnect_0_onchip_sram_s1_readdata),                   //                                                                .readdata
		.Onchip_SRAM_s1_writedata                                              (mm_interconnect_0_onchip_sram_s1_writedata),                  //                                                                .writedata
		.Onchip_SRAM_s1_byteenable                                             (mm_interconnect_0_onchip_sram_s1_byteenable),                 //                                                                .byteenable
		.Onchip_SRAM_s1_chipselect                                             (mm_interconnect_0_onchip_sram_s1_chipselect),                 //                                                                .chipselect
		.Onchip_SRAM_s1_clken                                                  (mm_interconnect_0_onchip_sram_s1_clken),                      //                                                                .clken
		.Onchip_SRAM_s2_address                                                (mm_interconnect_0_onchip_sram_s2_address),                    //                                                  Onchip_SRAM_s2.address
		.Onchip_SRAM_s2_write                                                  (mm_interconnect_0_onchip_sram_s2_write),                      //                                                                .write
		.Onchip_SRAM_s2_readdata                                               (mm_interconnect_0_onchip_sram_s2_readdata),                   //                                                                .readdata
		.Onchip_SRAM_s2_writedata                                              (mm_interconnect_0_onchip_sram_s2_writedata),                  //                                                                .writedata
		.Onchip_SRAM_s2_byteenable                                             (mm_interconnect_0_onchip_sram_s2_byteenable),                 //                                                                .byteenable
		.Onchip_SRAM_s2_chipselect                                             (mm_interconnect_0_onchip_sram_s2_chipselect),                 //                                                                .chipselect
		.Onchip_SRAM_s2_clken                                                  (mm_interconnect_0_onchip_sram_s2_clken),                      //                                                                .clken
		.SDRAM_s1_address                                                      (mm_interconnect_0_sdram_s1_address),                          //                                                        SDRAM_s1.address
		.SDRAM_s1_write                                                        (mm_interconnect_0_sdram_s1_write),                            //                                                                .write
		.SDRAM_s1_read                                                         (mm_interconnect_0_sdram_s1_read),                             //                                                                .read
		.SDRAM_s1_readdata                                                     (mm_interconnect_0_sdram_s1_readdata),                         //                                                                .readdata
		.SDRAM_s1_writedata                                                    (mm_interconnect_0_sdram_s1_writedata),                        //                                                                .writedata
		.SDRAM_s1_byteenable                                                   (mm_interconnect_0_sdram_s1_byteenable),                       //                                                                .byteenable
		.SDRAM_s1_readdatavalid                                                (mm_interconnect_0_sdram_s1_readdatavalid),                    //                                                                .readdatavalid
		.SDRAM_s1_waitrequest                                                  (mm_interconnect_0_sdram_s1_waitrequest),                      //                                                                .waitrequest
		.SDRAM_s1_chipselect                                                   (mm_interconnect_0_sdram_s1_chipselect),                       //                                                                .chipselect
		.vgasystem_0_char_buffer_slave_address                                 (mm_interconnect_0_vgasystem_0_char_buffer_slave_address),     //                                   vgasystem_0_char_buffer_slave.address
		.vgasystem_0_char_buffer_slave_write                                   (mm_interconnect_0_vgasystem_0_char_buffer_slave_write),       //                                                                .write
		.vgasystem_0_char_buffer_slave_read                                    (mm_interconnect_0_vgasystem_0_char_buffer_slave_read),        //                                                                .read
		.vgasystem_0_char_buffer_slave_readdata                                (mm_interconnect_0_vgasystem_0_char_buffer_slave_readdata),    //                                                                .readdata
		.vgasystem_0_char_buffer_slave_writedata                               (mm_interconnect_0_vgasystem_0_char_buffer_slave_writedata),   //                                                                .writedata
		.vgasystem_0_char_buffer_slave_byteenable                              (mm_interconnect_0_vgasystem_0_char_buffer_slave_byteenable),  //                                                                .byteenable
		.vgasystem_0_char_buffer_slave_waitrequest                             (mm_interconnect_0_vgasystem_0_char_buffer_slave_waitrequest), //                                                                .waitrequest
		.vgasystem_0_char_buffer_slave_chipselect                              (mm_interconnect_0_vgasystem_0_char_buffer_slave_chipselect)   //                                                                .chipselect
	);

	mysystem_mm_interconnect_1 mm_interconnect_1 (
		.arm_a9_hps_h2f_lw_axi_master_awid                                        (arm_a9_hps_h2f_lw_axi_master_awid),                                  //                                       arm_a9_hps_h2f_lw_axi_master.awid
		.arm_a9_hps_h2f_lw_axi_master_awaddr                                      (arm_a9_hps_h2f_lw_axi_master_awaddr),                                //                                                                   .awaddr
		.arm_a9_hps_h2f_lw_axi_master_awlen                                       (arm_a9_hps_h2f_lw_axi_master_awlen),                                 //                                                                   .awlen
		.arm_a9_hps_h2f_lw_axi_master_awsize                                      (arm_a9_hps_h2f_lw_axi_master_awsize),                                //                                                                   .awsize
		.arm_a9_hps_h2f_lw_axi_master_awburst                                     (arm_a9_hps_h2f_lw_axi_master_awburst),                               //                                                                   .awburst
		.arm_a9_hps_h2f_lw_axi_master_awlock                                      (arm_a9_hps_h2f_lw_axi_master_awlock),                                //                                                                   .awlock
		.arm_a9_hps_h2f_lw_axi_master_awcache                                     (arm_a9_hps_h2f_lw_axi_master_awcache),                               //                                                                   .awcache
		.arm_a9_hps_h2f_lw_axi_master_awprot                                      (arm_a9_hps_h2f_lw_axi_master_awprot),                                //                                                                   .awprot
		.arm_a9_hps_h2f_lw_axi_master_awvalid                                     (arm_a9_hps_h2f_lw_axi_master_awvalid),                               //                                                                   .awvalid
		.arm_a9_hps_h2f_lw_axi_master_awready                                     (arm_a9_hps_h2f_lw_axi_master_awready),                               //                                                                   .awready
		.arm_a9_hps_h2f_lw_axi_master_wid                                         (arm_a9_hps_h2f_lw_axi_master_wid),                                   //                                                                   .wid
		.arm_a9_hps_h2f_lw_axi_master_wdata                                       (arm_a9_hps_h2f_lw_axi_master_wdata),                                 //                                                                   .wdata
		.arm_a9_hps_h2f_lw_axi_master_wstrb                                       (arm_a9_hps_h2f_lw_axi_master_wstrb),                                 //                                                                   .wstrb
		.arm_a9_hps_h2f_lw_axi_master_wlast                                       (arm_a9_hps_h2f_lw_axi_master_wlast),                                 //                                                                   .wlast
		.arm_a9_hps_h2f_lw_axi_master_wvalid                                      (arm_a9_hps_h2f_lw_axi_master_wvalid),                                //                                                                   .wvalid
		.arm_a9_hps_h2f_lw_axi_master_wready                                      (arm_a9_hps_h2f_lw_axi_master_wready),                                //                                                                   .wready
		.arm_a9_hps_h2f_lw_axi_master_bid                                         (arm_a9_hps_h2f_lw_axi_master_bid),                                   //                                                                   .bid
		.arm_a9_hps_h2f_lw_axi_master_bresp                                       (arm_a9_hps_h2f_lw_axi_master_bresp),                                 //                                                                   .bresp
		.arm_a9_hps_h2f_lw_axi_master_bvalid                                      (arm_a9_hps_h2f_lw_axi_master_bvalid),                                //                                                                   .bvalid
		.arm_a9_hps_h2f_lw_axi_master_bready                                      (arm_a9_hps_h2f_lw_axi_master_bready),                                //                                                                   .bready
		.arm_a9_hps_h2f_lw_axi_master_arid                                        (arm_a9_hps_h2f_lw_axi_master_arid),                                  //                                                                   .arid
		.arm_a9_hps_h2f_lw_axi_master_araddr                                      (arm_a9_hps_h2f_lw_axi_master_araddr),                                //                                                                   .araddr
		.arm_a9_hps_h2f_lw_axi_master_arlen                                       (arm_a9_hps_h2f_lw_axi_master_arlen),                                 //                                                                   .arlen
		.arm_a9_hps_h2f_lw_axi_master_arsize                                      (arm_a9_hps_h2f_lw_axi_master_arsize),                                //                                                                   .arsize
		.arm_a9_hps_h2f_lw_axi_master_arburst                                     (arm_a9_hps_h2f_lw_axi_master_arburst),                               //                                                                   .arburst
		.arm_a9_hps_h2f_lw_axi_master_arlock                                      (arm_a9_hps_h2f_lw_axi_master_arlock),                                //                                                                   .arlock
		.arm_a9_hps_h2f_lw_axi_master_arcache                                     (arm_a9_hps_h2f_lw_axi_master_arcache),                               //                                                                   .arcache
		.arm_a9_hps_h2f_lw_axi_master_arprot                                      (arm_a9_hps_h2f_lw_axi_master_arprot),                                //                                                                   .arprot
		.arm_a9_hps_h2f_lw_axi_master_arvalid                                     (arm_a9_hps_h2f_lw_axi_master_arvalid),                               //                                                                   .arvalid
		.arm_a9_hps_h2f_lw_axi_master_arready                                     (arm_a9_hps_h2f_lw_axi_master_arready),                               //                                                                   .arready
		.arm_a9_hps_h2f_lw_axi_master_rid                                         (arm_a9_hps_h2f_lw_axi_master_rid),                                   //                                                                   .rid
		.arm_a9_hps_h2f_lw_axi_master_rdata                                       (arm_a9_hps_h2f_lw_axi_master_rdata),                                 //                                                                   .rdata
		.arm_a9_hps_h2f_lw_axi_master_rresp                                       (arm_a9_hps_h2f_lw_axi_master_rresp),                                 //                                                                   .rresp
		.arm_a9_hps_h2f_lw_axi_master_rlast                                       (arm_a9_hps_h2f_lw_axi_master_rlast),                                 //                                                                   .rlast
		.arm_a9_hps_h2f_lw_axi_master_rvalid                                      (arm_a9_hps_h2f_lw_axi_master_rvalid),                                //                                                                   .rvalid
		.arm_a9_hps_h2f_lw_axi_master_rready                                      (arm_a9_hps_h2f_lw_axi_master_rready),                                //                                                                   .rready
		.system_pll_sys_clk_clk                                                   (system_pll_sys_clk_clk),                                             //                                                 system_pll_sys_clk.clk
		.arm_a9_hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                                 // arm_a9_hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.jtag_uart_reset_reset_bridge_in_reset_reset                              (rst_controller_reset_out_reset),                                     //                              jtag_uart_reset_reset_bridge_in_reset.reset
		.vgasystem_0_sys_reset_reset_bridge_in_reset_reset                        (rst_controller_reset_out_reset),                                     //                        vgasystem_0_sys_reset_reset_bridge_in_reset.reset
		.jtag_uart_avalon_jtag_slave_address                                      (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),              //                                        jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                                        (mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),                //                                                                   .write
		.jtag_uart_avalon_jtag_slave_read                                         (mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),                 //                                                                   .read
		.jtag_uart_avalon_jtag_slave_readdata                                     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),             //                                                                   .readdata
		.jtag_uart_avalon_jtag_slave_writedata                                    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),            //                                                                   .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                                  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest),          //                                                                   .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                                   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),           //                                                                   .chipselect
		.vgasystem_0_char_buffer_control_slave_address                            (mm_interconnect_1_vgasystem_0_char_buffer_control_slave_address),    //                              vgasystem_0_char_buffer_control_slave.address
		.vgasystem_0_char_buffer_control_slave_write                              (mm_interconnect_1_vgasystem_0_char_buffer_control_slave_write),      //                                                                   .write
		.vgasystem_0_char_buffer_control_slave_read                               (mm_interconnect_1_vgasystem_0_char_buffer_control_slave_read),       //                                                                   .read
		.vgasystem_0_char_buffer_control_slave_readdata                           (mm_interconnect_1_vgasystem_0_char_buffer_control_slave_readdata),   //                                                                   .readdata
		.vgasystem_0_char_buffer_control_slave_writedata                          (mm_interconnect_1_vgasystem_0_char_buffer_control_slave_writedata),  //                                                                   .writedata
		.vgasystem_0_char_buffer_control_slave_byteenable                         (mm_interconnect_1_vgasystem_0_char_buffer_control_slave_byteenable), //                                                                   .byteenable
		.vgasystem_0_char_buffer_control_slave_chipselect                         (mm_interconnect_1_vgasystem_0_char_buffer_control_slave_chipselect), //                                                                   .chipselect
		.vgasystem_0_pixel_dma_control_slave_address                              (mm_interconnect_1_vgasystem_0_pixel_dma_control_slave_address),      //                                vgasystem_0_pixel_dma_control_slave.address
		.vgasystem_0_pixel_dma_control_slave_write                                (mm_interconnect_1_vgasystem_0_pixel_dma_control_slave_write),        //                                                                   .write
		.vgasystem_0_pixel_dma_control_slave_read                                 (mm_interconnect_1_vgasystem_0_pixel_dma_control_slave_read),         //                                                                   .read
		.vgasystem_0_pixel_dma_control_slave_readdata                             (mm_interconnect_1_vgasystem_0_pixel_dma_control_slave_readdata),     //                                                                   .readdata
		.vgasystem_0_pixel_dma_control_slave_writedata                            (mm_interconnect_1_vgasystem_0_pixel_dma_control_slave_writedata),    //                                                                   .writedata
		.vgasystem_0_pixel_dma_control_slave_byteenable                           (mm_interconnect_1_vgasystem_0_pixel_dma_control_slave_byteenable)    //                                                                   .byteenable
	);

	mysystem_irq_mapper irq_mapper (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.sender_irq    (arm_a9_hps_f2h_irq0_irq)   //    sender.irq
	);

	mysystem_irq_mapper_001 irq_mapper_001 (
		.clk        (),                        //       clk.clk
		.reset      (),                        // clk_reset.reset
		.sender_irq (arm_a9_hps_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (system_pll_reset_source_reset),      // reset_in0.reset
		.reset_in1      (~arm_a9_hps_h2f_reset_reset),        // reset_in1.reset
		.clk            (system_pll_sys_clk_clk),             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (system_pll_reset_source_reset),      // reset_in0.reset
		.reset_in1      (~arm_a9_hps_h2f_reset_reset),        // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.clk            (system_pll_sys_clk_clk),             //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
